module xor_tb;
    reg a, b;
    wire y;

    xorgate dut (
        .a(a),
        .b(b),
        .y(y)
    );

    initial begin
        $dumpfile("xor_wave.vcd");
        $dumpvars(0, xor_tb);

        a = 0;
        b = 0;
        #10;
        a = 0;
        b = 1;
        #10;
        a = 1;
        b = 0;
        #10;
        a = 1;
        b = 1;
        #10;
        $finish;
    end
endmodule
