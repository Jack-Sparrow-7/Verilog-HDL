module nand_gate(
    a,b,y
);

input a,b;
output y;

nand(y,a,b);
    
endmodule