module nor_gate(a,b,y);
    input a,b;
    output y;

    nor object(y,a,b);

endmodule


